module signExtend
(	input signed [15:0] in,
	output signed [31:0] out
	);

assign out = in;

endmodule: signExtend